`define WB_ADDR_I 4
`define WB_DAT_I 8
`define WB_DAT_O 8
